module tb_adder_16x23bit;
    reg [22:0] in [15:0];
    wire [22:0] sum;
    wire carry_out;

    adder_16x23bit uut (
        .in(in),
        .sum(sum),
        .carry_out(carry_out)
    );

    initial begin
        $monitor("Time = %0d, sum = %023b, carry_out = %b", $time, sum, carry_out);

        // Test case: all zeros
        in[0] = 23'b00000000000000000000000; 
        in[1] = 23'b00000000000000000000000; 
        in[2] = 23'b00000000000000000000000; 
        in[3] = 23'b00000000000000000000000; 
        in[4] = 23'b00000000000000000000000; 
        in[5] = 23'b00000000000000000000000; 
        in[6] = 23'b00000000000000000000000; 
        in[7] = 23'b00000000000000000000000; 
        in[8] = 23'b00000000000000000000000; 
        in[9] = 23'b00000000000000000000000; 
        in[10] = 23'b00000000000000000000000; 
        in[11] = 23'b00000000000000000000000; 
        in[12] = 23'b00000000000000000000000; 
        in[13] = 23'b00000000000000000000000; 
        in[14] = 23'b00000000000000000000000; 
        in[15] = 23'b00000000000000000000000; 
        #10;

        // Test case: all ones
        in[0] = 23'b00000000000000000000001; 
        in[1] = 23'b00000000000000000000001; 
        in[2] = 23'b00000000000000000000001; 
        in[3] = 23'b00000000000000000000001; 
        in[4] = 23'b00000000000000000000001; 
        in[5] = 23'b00000000000000000000001; 
        in[6] = 23'b00000000000000000000001; 
        in[7] = 23'b00000000000000000000001; 
        in[8] = 23'b00000000000000000000001; 
        in[9] = 23'b00000000000000000000001; 
        in[10] = 23'b00000000000000000000001; 
        in[11] = 23'b00000000000000000000001; 
        in[12] = 23'b00000000000000000000001; 
        in[13] = 23'b00000000000000000000001; 
        in[14] = 23'b00000000000000000000001; 
        in[15] = 23'b00000000000000000000001; 
        #10;

        // Test case: random values
        in[0] = 23'b10101010101010101010101; 
        in[1] = 23'b01010101010101010101010; 
        in[2] = 23'b11100011100011100011100; 
        in[3] = 23'b00011100011100011100011; 
        in[4] = 23'b10010010010010010010010; 
        in[5] = 23'b01101101101101101101101; 
        in[6] = 23'b00000000000000000000000; 
        in[7] = 23'b11111111111111111111111; 
        in[8] = 23'b00100100100100100100100; 
        in[9] = 23'b01001001001001001001001; 
        in[10] = 23'b11111111111111111111111; 
        in[11] = 23'b00000000000000000000000; 
        in[12] = 23'b10101010101010101010101; 
        in[13] = 23'b01010101010101010101010; 
        in[14] = 23'b11100011100011100011100; 
        in[15] = 23'b00011100011100011100011; 
        #10;

        $finish;
    end
endmodule
