module tb_adder_23bit;
    reg [22:0] a;
    reg [22:0] b;
    wire [22:0] sum;
    wire carry_out;

    adder_23bit uut (
        .a(a),
        .b(b),
        .sum(sum),
        .carry_out(carry_out)
    );

    initial begin
        $monitor("Time = %0d, a = %023b, b = %023b, sum = %023b, carry_out = %b", $time, a, b, sum, carry_out);

        // Test cases with two's complement signed numbers
        a = 23'b00000000000000000000001; b = 23'b00000000000000000000001; #10;
        a = 23'b11111111111111111111111; b = 23'b00000000000000000000001; #10;
        a = 23'b10101010101010101010101; b = 23'b01010101010101010101010; #10;
        a = 23'b11111111111111111111111; b = 23'b11111111111111111111111; #10;

        // Test negative numbers (in two's complement)
        a = 23'b11111111111111111111110; b = 23'b00000000000000000000001; #10; // -2 + 1
        a = 23'b11111111111111111110000; b = 23'b00000000000000000001000; #10; // -16 + 8

        // Test carry out
        a = 23'b01111111111111111111111; b = 23'b00000000000000000000001; #10; // 4194303 + 1

        // Test overflow
        a = 23'b01111111111111111111111; b = 23'b01111111111111111111111; #10; // 4194303 + 4194303

        // Test all zeros
        a = 23'b00000000000000000000000; b = 23'b00000000000000000000000; #10;

        // Test random values
        a = 23'b01010101010101010101010; b = 23'b00101010101010101010101; #10;
        a = 23'b11100011100011100011100; b = 23'b00011100011100011100011; #10;

        $finish;
    end
endmodule
